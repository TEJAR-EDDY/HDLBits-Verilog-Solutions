module top_module ( 
    input clk, 
    input [7:0] d, 
    input [1:0] sel, 
    output [7:0] q 
);
 wire [7:0] q1, q2, q3;  // Wires to connect between DFF stages

    // Instantiate three 8-bit D flip-flop modules
    my_dff8 dff1 ( .clk(clk), .d(d),   .q(q1) );
    my_dff8 dff2 ( .clk(clk), .d(q1),  .q(q2) );
    my_dff8 dff3 ( .clk(clk), .d(q2),  .q(q3) );

    // 4-to-1 multiplexer to select output based on sel
    always @(*) begin
        case (sel)
            2'b00: q = d;   // No delay
            2'b01: q = q1;  // 1-cycle delay
            2'b10: q = q2;  // 2-cycle delay
            2'b11: q = q3;  // 3-cycle delay
        endcase
    end

endmodule
